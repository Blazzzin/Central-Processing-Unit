library verilog;
use verilog.vl_types.all;
entity problem2_vlg_vec_tst is
end problem2_vlg_vec_tst;
