library verilog;
use verilog.vl_types.all;
entity problem1_vlg_vec_tst is
end problem1_vlg_vec_tst;
