library verilog;
use verilog.vl_types.all;
entity ALU1_vlg_vec_tst is
end ALU1_vlg_vec_tst;
